// test to verify assign statements

module testmodule(x1,x2,x3,x4,y1,y2,y3,y4);

input x1;
input x2;
input x3;
input x4;
output y1;
output y2;
output y3;
output y4;

assign y1 = x1;
assign y2 = x2;
assign y3 = x3;
assign y4 = x4;

endmodule
