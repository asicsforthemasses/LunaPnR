# SPDX-FileCopyrightText: 2021-2025 Niels Moseley <asicsforthemasses@gmail.com>
#
# SPDX-License-Identifier: GPL-3.0-only
#

VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS

USEMINSPACING OBS ON ;
USEMINSPACING PIN OFF ;
CLEARANCEMEASURE EUCLIDEAN ;

MANUFACTURINGGRID 0.05 ;

SITE  core
    CLASS	CORE ;
    SYMMETRY	Y ;
    SIZE	0.800 BY 10.000 ;
END  core

MACRO TIEHI
  CLASS  CORE ;
  FOREIGN INVX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.600 BY 10.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.200 -0.300 0.600 1.600 ;
        RECT -0.200 -0.300 1.800 0.300 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 1.000 0.600 1.400 9.400 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.200 7.400 0.600 10.300 ;
        RECT -0.200 9.700 1.800 10.300 ;
    END
  END vdd
END TIEHI

MACRO TIELO
  CLASS  CORE ;
  FOREIGN INVX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.600 BY 10.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.200 -0.300 0.600 1.600 ;
        RECT -0.200 -0.300 1.800 0.300 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 1.000 0.600 1.400 9.400 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.200 7.400 0.600 10.300 ;
        RECT -0.200 9.700 1.800 10.300 ;
    END
  END vdd
END TIELO

MACRO __PIN
  CLASS  CORE ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.00 BY 4.00 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN Y
    DIRECTION INOUT ;
    PORT
      LAYER metal1 ;
        RECT 1.000 1.000 3.00 3.00 ;
    END
  END Y
END __PIN

END LIBRARY
