# SPDX-FileCopyrightText: 2021-2025 Niels Moseley <asicsforthemasses@gmail.com>
#
# SPDX-License-Identifier: GPL-3.0-only
#

VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS

USEMINSPACING OBS ON ;
USEMINSPACING PIN OFF ;
CLEARANCEMEASURE EUCLIDEAN ;

MANUFACTURINGGRID 0.05 ;

SITE  core
    CLASS	CORE ;
    SYMMETRY	Y ;
    SIZE	0.800 BY 10.000 ;
END  core

MACRO PADNC5
  CLASS  PAD ;
  FOREIGN PADNC5 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 300.000 ;
  SYMMETRY R90 ;
  SITE IO ;
  OBS
      LAYER metal4 ;
        RECT 0.600 0.600 4.400 299.400 ;
      LAYER metal3 ;
        RECT 0.600 0.600 4.400 299.400 ;
      LAYER metal2 ;
        RECT 0.000 0.000 5.000 72.400 ;
        RECT 0.000 76.800 5.000 97.800 ;
        RECT 0.000 104.200 5.000 125.200 ;
        RECT 0.000 129.600 5.000 202.000 ;
        RECT 0.600 0.000 4.400 299.400 ;
      LAYER metal1 ;
        RECT 0.000 0.000 5.000 97.800 ;
        RECT 0.000 104.200 5.000 202.000 ;
        RECT 0.600 0.000 4.400 299.400 ;
  END
END PADNC5

MACRO PADNC10
  CLASS  PAD ;
  FOREIGN PADNC10 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 300.000 ;
  SYMMETRY R90 ;
  SITE IO ;
  OBS
      LAYER metal4 ;
        RECT 0.600 0.600 9.400 299.400 ;
      LAYER metal3 ;
        RECT 0.600 0.600 9.400 299.400 ;
      LAYER metal2 ;
        RECT 0.000 0.000 10.000 72.400 ;
        RECT 0.000 76.800 10.000 97.800 ;
        RECT 0.000 104.200 10.000 125.200 ;
        RECT 0.000 129.600 10.000 202.000 ;
        RECT 0.600 0.000 9.400 299.400 ;
      LAYER metal1 ;
        RECT 0.000 0.000 10.000 97.800 ;
        RECT 0.000 104.200 10.000 202.000 ;
        RECT 0.600 0.000 9.400 299.400 ;
  END
END PADNC10

MACRO PADNC50
  CLASS  PAD ;
  FOREIGN PADNC50 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 50.000 BY 300.000 ;
  SYMMETRY R90 ;
  SITE IO ;
  OBS
      LAYER metal4 ;
        RECT 0.600 0.600 49.400 299.400 ;
      LAYER metal3 ;
        RECT 0.600 0.600 49.400 299.400 ;
      LAYER metal2 ;
        RECT 0.000 0.000 50.000 72.400 ;
        RECT 0.000 76.800 50.000 97.800 ;
        RECT 0.000 104.200 50.000 125.200 ;
        RECT 0.000 129.600 50.000 202.000 ;
        RECT 0.600 0.000 49.400 299.400 ;
      LAYER metal1 ;
        RECT 0.000 0.000 50.000 97.800 ;
        RECT 0.000 104.200 50.000 202.000 ;
        RECT 0.600 0.000 49.400 299.400 ;
  END
END PADNC50

END LIBRARY
